module simpleor(f,x,y);
    input x,y;
    output f;
    or a1(f,x,y);
endmodule
