module simpleand(f,x,y);
    input x,y;
    output f;
    and a1(f,x,y);
endmodule
