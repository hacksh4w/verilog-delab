module gray2bin_tb();

reg g3,g2,g1,g0;
wire b3,b2,b1,b0;

gray2bin dut(g3,g2,g1,g0,b3,b2,b1,b0);

initial
    begin
        g3 = 0; g2 = 0; g1 = 0; g0 = 0; #20
        g3 = 0; g2 = 0; g1 = 0; g0 = 1; #20
        g3 = 0; g2 = 0; g1 = 1; g0 = 0; #20
        g3 = 0; g2 = 0; g1 = 1; g0 = 1; #20
        g3 = 0; g2 = 1; g1 = 0; g0 = 0; #20
        g3 = 0; g2 = 1; g1 = 0; g0 = 1; #20
        g3 = 0; g2 = 1; g1 = 1; g0 = 0; #20
        g3 = 0; g2 = 1; g1 = 1; g0 = 1; #20
        g3 = 1; g2 = 0; g1 = 0; g0 = 0; #20
        g3 = 1; g2 = 0; g1 = 0; g0 = 1; #20
        g3 = 1; g2 = 0; g1 = 1; g0 = 0; #20
        g3 = 1; g2 = 0; g1 = 1; g0 = 1; #20
        g3 = 1; g2 = 1; g1 = 0; g0 = 0; #20
        g3 = 1; g2 = 1; g1 = 0; g0 = 1; #20
        g3 = 1; g2 = 1; g1 = 1; g0 = 0; #20
        g3 = 1; g2 = 1; g1 = 1; g0 = 1; #20
        $finish(); 
    end
endmodule
