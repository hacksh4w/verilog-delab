module nand_s(a,b,z);
input a,b;
output z;

nand a1(z,a,b);
                
endmodule
