module xnor_s(a,b,y);
input a,b;
output y;

xnor b1(y,a,b);
                
endmodule
