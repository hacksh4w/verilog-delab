module not_gate_s(a,y);
input a;
output y;

not a1(y,a);         
endmodule
