module bin2gray_tb();

reg b0,b1,b2,b3;
wire g0,g1,g2,g3;

bin2gray dut(b3,b2,b1,b0,g3,g2,g1,g0);

initial
    begin
        b3 = 0; b2 = 0; b1 = 0; b0 = 0; #20
        b3 = 0; b2 = 0; b1 = 0; b0 = 1; #20
        b3 = 0; b2 = 0; b1 = 1; b0 = 0; #20
        b3 = 0; b2 = 0; b1 = 1; b0 = 1; #20
        b3 = 0; b2 = 1; b1 = 0; b0 = 0; #20
        b3 = 0; b2 = 1; b1 = 0; b0 = 1; #20
        b3 = 0; b2 = 1; b1 = 1; b0 = 0; #20
        b3 = 0; b2 = 1; b1 = 1; b0 = 1; #20
        b3 = 1; b2 = 0; b1 = 0; b0 = 0; #20
        b3 = 1; b2 = 0; b1 = 0; b0 = 1; #20
        b3 = 1; b2 = 0; b1 = 1; b0 = 0; #20
        b3 = 1; b2 = 0; b1 = 1; b0 = 1; #20
        b3 = 1; b2 = 1; b1 = 0; b0 = 0; #20
        b3 = 1; b2 = 1; b1 = 0; b0 = 1; #20
        b3 = 1; b2 = 1; b1 = 1; b0 = 0; #20
        b3 = 1; b2 = 1; b1 = 1; b0 = 1; #20
        $finish(); 
    end
endmodule
